`timescale 1ns / 1ns
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05.12.2024 14:02:24
// Design Name: 
// Module Name: FeederTest
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module FeederTest(

    );
    
    reg [7:0] character_id;
    wire [3:0] row;
    wire [5:0] col;
    wire push_up;
    wire reset_call;
    reg clock;
    
    CharacterFeeder characterFeeder(row,col,character_id,push_up,reset_call,1,clock);
    
    initial begin
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
        #1 clock = 0;
        #1 clock = 1;
    end
    
endmodule
