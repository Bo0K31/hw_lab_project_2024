`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 27.11.2024 09:13:01
// Design Name: 
// Module Name: ChracterPlaneTest
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ChracterPlaneTest(

    );
    wire [3:0] row;
    wire [5:0] column;
    wire [7:0] character_id;
    reg [3:0] _row;
    reg [5:0] _column;
    reg [7:0] _character_id;
    reg reset;
    reg clock;
    reg we;
    
    reg [3:0] a;
    reg [5:0] b;
    reg [7:0] c;
    
    CharacterPlane characterPlane(character_id,row,column,_character_id,_row,_column,we,reset,clock);
    
    assign row = a;
    assign column = b;
    always@(row, column, character_id) begin
        c <= character_id;
    end
    
    initial begin
        we = 0; _row = 0; _column = 0; reset = 0; clock = 0;
        #10; we = 1; _row = 0; _column = 0; _character_id = 1;
        #1; clock = 1;
        #1; clock = 0;
        #10; we = 1; _row = 0; _column = 1; _character_id = 2;
        #1; clock = 1;
        #1; clock = 0;
        #10; we = 1; _row = 0; _column = 2; _character_id = 3;
        #1; clock = 1;
        #1; clock = 0;
        #10; we = 1; _row = 0; _column = 3; _character_id = 4;
        #1; clock = 1;
        #1; clock = 0;
        #1; a = 0; b = 0;
        
        #10; reset = 1; we= 0;
        
#1; a = 0; b = 1;
#1; a = 0; b = 2;
#1; a = 0; b = 3;
#1; a = 0; b = 4;
#1; a = 0; b = 5;
#1; a = 0; b = 6;
#1; a = 0; b = 7;
#1; a = 0; b = 8;
#1; a = 0; b = 9;
#1; a = 0; b = 10;
#1; a = 0; b = 11;
#1; a = 0; b = 12;
#1; a = 0; b = 13;
#1; a = 0; b = 14;
#1; a = 0; b = 15;
#1; a = 0; b = 16;
#1; a = 0; b = 17;
#1; a = 0; b = 18;
#1; a = 0; b = 19;
#1; a = 0; b = 20;
#1; a = 0; b = 21;
#1; a = 0; b = 22;
#1; a = 0; b = 23;
#1; a = 0; b = 24;
#1; a = 0; b = 25;
#1; a = 0; b = 26;
#1; a = 0; b = 27;
#1; a = 0; b = 28;
#1; a = 0; b = 29;
#1; a = 0; b = 30;
#1; a = 0; b = 31;
#1; a = 0; b = 32;
#1; a = 0; b = 33;
#1; a = 0; b = 34;
#1; a = 0; b = 35;
#1; a = 0; b = 36;
#1; a = 0; b = 37;
#1; a = 0; b = 38;
#1; a = 0; b = 39;
#1; a = 1; b = 0;
#1; a = 1; b = 1;
#1; a = 1; b = 2;
#1; a = 1; b = 3;
#1; a = 1; b = 4;
#1; a = 1; b = 5;
#1; a = 1; b = 6;
#1; a = 1; b = 7;
#1; a = 1; b = 8;
#1; a = 1; b = 9;
#1; a = 1; b = 10;
#1; a = 1; b = 11;
#1; a = 1; b = 12;
#1; a = 1; b = 13;
#1; a = 1; b = 14;
#1; a = 1; b = 15;
#1; a = 1; b = 16;
#1; a = 1; b = 17;
#1; a = 1; b = 18;
#1; a = 1; b = 19;
#1; a = 1; b = 20;
#1; a = 1; b = 21;
#1; a = 1; b = 22;
#1; a = 1; b = 23;
#1; a = 1; b = 24;
#1; a = 1; b = 25;
#1; a = 1; b = 26;
#1; a = 1; b = 27;
#1; a = 1; b = 28;
#1; a = 1; b = 29;
#1; a = 1; b = 30;
#1; a = 1; b = 31;
#1; a = 1; b = 32;
#1; a = 1; b = 33;
#1; a = 1; b = 34;
#1; a = 1; b = 35;
#1; a = 1; b = 36;
#1; a = 1; b = 37;
#1; a = 1; b = 38;
#1; a = 1; b = 39;
#1; a = 2; b = 0;
#1; a = 2; b = 1;
#1; a = 2; b = 2;
#1; a = 2; b = 3;
#1; a = 2; b = 4;
#1; a = 2; b = 5;
#1; a = 2; b = 6;
#1; a = 2; b = 7;
#1; a = 2; b = 8;
#1; a = 2; b = 9;
#1; a = 2; b = 10;
#1; a = 2; b = 11;
#1; a = 2; b = 12;
#1; a = 2; b = 13;
#1; a = 2; b = 14;
#1; a = 2; b = 15;
#1; a = 2; b = 16;
#1; a = 2; b = 17;
#1; a = 2; b = 18;
#1; a = 2; b = 19;
#1; a = 2; b = 20;
#1; a = 2; b = 21;
#1; a = 2; b = 22;
#1; a = 2; b = 23;
#1; a = 2; b = 24;
#1; a = 2; b = 25;
#1; a = 2; b = 26;
#1; a = 2; b = 27;
#1; a = 2; b = 28;
#1; a = 2; b = 29;
#1; a = 2; b = 30;
#1; a = 2; b = 31;
#1; a = 2; b = 32;
#1; a = 2; b = 33;
#1; a = 2; b = 34;
#1; a = 2; b = 35;
#1; a = 2; b = 36;
#1; a = 2; b = 37;
#1; a = 2; b = 38;
#1; a = 2; b = 39;
#1; a = 3; b = 0;
#1; a = 3; b = 1;
#1; a = 3; b = 2;
#1; a = 3; b = 3;
#1; a = 3; b = 4;
#1; a = 3; b = 5;
#1; a = 3; b = 6;
#1; a = 3; b = 7;
#1; a = 3; b = 8;
#1; a = 3; b = 9;
#1; a = 3; b = 10;
#1; a = 3; b = 11;
#1; a = 3; b = 12;
#1; a = 3; b = 13;
#1; a = 3; b = 14;
#1; a = 3; b = 15;
#1; a = 3; b = 16;
#1; a = 3; b = 17;
#1; a = 3; b = 18;
#1; a = 3; b = 19;
#1; a = 3; b = 20;
#1; a = 3; b = 21;
#1; a = 3; b = 22;
#1; a = 3; b = 23;
#1; a = 3; b = 24;
#1; a = 3; b = 25;
#1; a = 3; b = 26;
#1; a = 3; b = 27;
#1; a = 3; b = 28;
#1; a = 3; b = 29;
#1; a = 3; b = 30;
#1; a = 3; b = 31;
#1; a = 3; b = 32;
#1; a = 3; b = 33;
#1; a = 3; b = 34;
#1; a = 3; b = 35;
#1; a = 3; b = 36;
#1; a = 3; b = 37;
#1; a = 3; b = 38;
#1; a = 3; b = 39;
#1; a = 4; b = 0;
#1; a = 4; b = 1;
#1; a = 4; b = 2;
#1; a = 4; b = 3;
#1; a = 4; b = 4;
#1; a = 4; b = 5;
#1; a = 4; b = 6;
#1; a = 4; b = 7;
#1; a = 4; b = 8;
#1; a = 4; b = 9;
#1; a = 4; b = 10;
#1; a = 4; b = 11;
#1; a = 4; b = 12;
#1; a = 4; b = 13;
#1; a = 4; b = 14;
#1; a = 4; b = 15;
#1; a = 4; b = 16;
#1; a = 4; b = 17;
#1; a = 4; b = 18;
#1; a = 4; b = 19;
#1; a = 4; b = 20;
#1; a = 4; b = 21;
#1; a = 4; b = 22;
#1; a = 4; b = 23;
#1; a = 4; b = 24;
#1; a = 4; b = 25;
#1; a = 4; b = 26;
#1; a = 4; b = 27;
#1; a = 4; b = 28;
#1; a = 4; b = 29;
#1; a = 4; b = 30;
#1; a = 4; b = 31;
#1; a = 4; b = 32;
#1; a = 4; b = 33;
#1; a = 4; b = 34;
#1; a = 4; b = 35;
#1; a = 4; b = 36;
#1; a = 4; b = 37;
#1; a = 4; b = 38;
#1; a = 4; b = 39;
#1; a = 5; b = 0;
#1; a = 5; b = 1;
#1; a = 5; b = 2;
#1; a = 5; b = 3;
#1; a = 5; b = 4;
#1; a = 5; b = 5;
#1; a = 5; b = 6;
#1; a = 5; b = 7;
#1; a = 5; b = 8;
#1; a = 5; b = 9;
#1; a = 5; b = 10;
#1; a = 5; b = 11;
#1; a = 5; b = 12;
#1; a = 5; b = 13;
#1; a = 5; b = 14;
#1; a = 5; b = 15;
#1; a = 5; b = 16;
#1; a = 5; b = 17;
#1; a = 5; b = 18;
#1; a = 5; b = 19;
#1; a = 5; b = 20;
#1; a = 5; b = 21;
#1; a = 5; b = 22;
#1; a = 5; b = 23;
#1; a = 5; b = 24;
#1; a = 5; b = 25;
#1; a = 5; b = 26;
#1; a = 5; b = 27;
#1; a = 5; b = 28;
#1; a = 5; b = 29;
#1; a = 5; b = 30;
#1; a = 5; b = 31;
#1; a = 5; b = 32;
#1; a = 5; b = 33;
#1; a = 5; b = 34;
#1; a = 5; b = 35;
#1; a = 5; b = 36;
#1; a = 5; b = 37;
#1; a = 5; b = 38;
#1; a = 5; b = 39;
#1; a = 6; b = 0;
#1; a = 6; b = 1;
#1; a = 6; b = 2;
#1; a = 6; b = 3;
#1; a = 6; b = 4;
#1; a = 6; b = 5;
#1; a = 6; b = 6;
#1; a = 6; b = 7;
#1; a = 6; b = 8;
#1; a = 6; b = 9;
#1; a = 6; b = 10;
#1; a = 6; b = 11;
#1; a = 6; b = 12;
#1; a = 6; b = 13;
#1; a = 6; b = 14;
#1; a = 6; b = 15;
#1; a = 6; b = 16;
#1; a = 6; b = 17;
#1; a = 6; b = 18;
#1; a = 6; b = 19;
#1; a = 6; b = 20;
#1; a = 6; b = 21;
#1; a = 6; b = 22;
#1; a = 6; b = 23;
#1; a = 6; b = 24;
#1; a = 6; b = 25;
#1; a = 6; b = 26;
#1; a = 6; b = 27;
#1; a = 6; b = 28;
#1; a = 6; b = 29;
#1; a = 6; b = 30;
#1; a = 6; b = 31;
#1; a = 6; b = 32;
#1; a = 6; b = 33;
#1; a = 6; b = 34;
#1; a = 6; b = 35;
#1; a = 6; b = 36;
#1; a = 6; b = 37;
#1; a = 6; b = 38;
#1; a = 6; b = 39;
#1; a = 7; b = 0;
#1; a = 7; b = 1;
#1; a = 7; b = 2;
#1; a = 7; b = 3;
#1; a = 7; b = 4;
#1; a = 7; b = 5;
#1; a = 7; b = 6;
#1; a = 7; b = 7;
#1; a = 7; b = 8;
#1; a = 7; b = 9;
#1; a = 7; b = 10;
#1; a = 7; b = 11;
#1; a = 7; b = 12;
#1; a = 7; b = 13;
#1; a = 7; b = 14;
#1; a = 7; b = 15;
#1; a = 7; b = 16;
#1; a = 7; b = 17;
#1; a = 7; b = 18;
#1; a = 7; b = 19;
#1; a = 7; b = 20;
#1; a = 7; b = 21;
#1; a = 7; b = 22;
#1; a = 7; b = 23;
#1; a = 7; b = 24;
#1; a = 7; b = 25;
#1; a = 7; b = 26;
#1; a = 7; b = 27;
#1; a = 7; b = 28;
#1; a = 7; b = 29;
#1; a = 7; b = 30;
#1; a = 7; b = 31;
#1; a = 7; b = 32;
#1; a = 7; b = 33;
#1; a = 7; b = 34;
#1; a = 7; b = 35;
#1; a = 7; b = 36;
#1; a = 7; b = 37;
#1; a = 7; b = 38;
#1; a = 7; b = 39;
#1; a = 8; b = 0;
#1; a = 8; b = 1;
#1; a = 8; b = 2;
#1; a = 8; b = 3;
#1; a = 8; b = 4;
#1; a = 8; b = 5;
#1; a = 8; b = 6;
#1; a = 8; b = 7;
#1; a = 8; b = 8;
#1; a = 8; b = 9;
#1; a = 8; b = 10;
#1; a = 8; b = 11;
#1; a = 8; b = 12;
#1; a = 8; b = 13;
#1; a = 8; b = 14;
#1; a = 8; b = 15;
#1; a = 8; b = 16;
#1; a = 8; b = 17;
#1; a = 8; b = 18;
#1; a = 8; b = 19;
#1; a = 8; b = 20;
#1; a = 8; b = 21;
#1; a = 8; b = 22;
#1; a = 8; b = 23;
#1; a = 8; b = 24;
#1; a = 8; b = 25;
#1; a = 8; b = 26;
#1; a = 8; b = 27;
#1; a = 8; b = 28;
#1; a = 8; b = 29;
#1; a = 8; b = 30;
#1; a = 8; b = 31;
#1; a = 8; b = 32;
#1; a = 8; b = 33;
#1; a = 8; b = 34;
#1; a = 8; b = 35;
#1; a = 8; b = 36;
#1; a = 8; b = 37;
#1; a = 8; b = 38;
#1; a = 8; b = 39;
#1; a = 9; b = 0;
#1; a = 9; b = 1;
#1; a = 9; b = 2;
#1; a = 9; b = 3;
#1; a = 9; b = 4;
#1; a = 9; b = 5;
#1; a = 9; b = 6;
#1; a = 9; b = 7;
#1; a = 9; b = 8;
#1; a = 9; b = 9;
#1; a = 9; b = 10;
#1; a = 9; b = 11;
#1; a = 9; b = 12;
#1; a = 9; b = 13;
#1; a = 9; b = 14;
#1; a = 9; b = 15;
#1; a = 9; b = 16;
#1; a = 9; b = 17;
#1; a = 9; b = 18;
#1; a = 9; b = 19;
#1; a = 9; b = 20;
#1; a = 9; b = 21;
#1; a = 9; b = 22;
#1; a = 9; b = 23;
#1; a = 9; b = 24;
#1; a = 9; b = 25;
#1; a = 9; b = 26;
#1; a = 9; b = 27;
#1; a = 9; b = 28;
#1; a = 9; b = 29;
#1; a = 9; b = 30;
#1; a = 9; b = 31;
#1; a = 9; b = 32;
#1; a = 9; b = 33;
#1; a = 9; b = 34;
#1; a = 9; b = 35;
#1; a = 9; b = 36;
#1; a = 9; b = 37;
#1; a = 9; b = 38;
#1; a = 9; b = 39;
#1; a = 10; b = 0;
#1; a = 10; b = 1;
#1; a = 10; b = 2;
#1; a = 10; b = 3;
#1; a = 10; b = 4;
#1; a = 10; b = 5;
#1; a = 10; b = 6;
#1; a = 10; b = 7;
#1; a = 10; b = 8;
#1; a = 10; b = 9;
#1; a = 10; b = 10;
#1; a = 10; b = 11;
#1; a = 10; b = 12;
#1; a = 10; b = 13;
#1; a = 10; b = 14;
#1; a = 10; b = 15;
#1; a = 10; b = 16;
#1; a = 10; b = 17;
#1; a = 10; b = 18;
#1; a = 10; b = 19;
#1; a = 10; b = 20;
#1; a = 10; b = 21;
#1; a = 10; b = 22;
#1; a = 10; b = 23;
#1; a = 10; b = 24;
#1; a = 10; b = 25;
#1; a = 10; b = 26;
#1; a = 10; b = 27;
#1; a = 10; b = 28;
#1; a = 10; b = 29;
#1; a = 10; b = 30;
#1; a = 10; b = 31;
#1; a = 10; b = 32;
#1; a = 10; b = 33;
#1; a = 10; b = 34;
#1; a = 10; b = 35;
#1; a = 10; b = 36;
#1; a = 10; b = 37;
#1; a = 10; b = 38;
#1; a = 10; b = 39;
#1; a = 11; b = 0;
#1; a = 11; b = 1;
#1; a = 11; b = 2;
#1; a = 11; b = 3;
#1; a = 11; b = 4;
#1; a = 11; b = 5;
#1; a = 11; b = 6;
#1; a = 11; b = 7;
#1; a = 11; b = 8;
#1; a = 11; b = 9;
#1; a = 11; b = 10;
#1; a = 11; b = 11;
#1; a = 11; b = 12;
#1; a = 11; b = 13;
#1; a = 11; b = 14;
#1; a = 11; b = 15;
#1; a = 11; b = 16;
#1; a = 11; b = 17;
#1; a = 11; b = 18;
#1; a = 11; b = 19;
#1; a = 11; b = 20;
#1; a = 11; b = 21;
#1; a = 11; b = 22;
#1; a = 11; b = 23;
#1; a = 11; b = 24;
#1; a = 11; b = 25;
#1; a = 11; b = 26;
#1; a = 11; b = 27;
#1; a = 11; b = 28;
#1; a = 11; b = 29;
#1; a = 11; b = 30;
#1; a = 11; b = 31;
#1; a = 11; b = 32;
#1; a = 11; b = 33;
#1; a = 11; b = 34;
#1; a = 11; b = 35;
#1; a = 11; b = 36;
#1; a = 11; b = 37;
#1; a = 11; b = 38;
#1; a = 11; b = 39;
#1; a = 12; b = 0;
#1; a = 12; b = 1;
#1; a = 12; b = 2;
#1; a = 12; b = 3;
#1; a = 12; b = 4;
#1; a = 12; b = 5;
#1; a = 12; b = 6;
#1; a = 12; b = 7;
#1; a = 12; b = 8;
#1; a = 12; b = 9;
#1; a = 12; b = 10;
#1; a = 12; b = 11;
#1; a = 12; b = 12;
#1; a = 12; b = 13;
#1; a = 12; b = 14;
#1; a = 12; b = 15;
#1; a = 12; b = 16;
#1; a = 12; b = 17;
#1; a = 12; b = 18;
#1; a = 12; b = 19;
#1; a = 12; b = 20;
#1; a = 12; b = 21;
#1; a = 12; b = 22;
#1; a = 12; b = 23;
#1; a = 12; b = 24;
#1; a = 12; b = 25;
#1; a = 12; b = 26;
#1; a = 12; b = 27;
#1; a = 12; b = 28;
#1; a = 12; b = 29;
#1; a = 12; b = 30;
#1; a = 12; b = 31;
#1; a = 12; b = 32;
#1; a = 12; b = 33;
#1; a = 12; b = 34;
#1; a = 12; b = 35;
#1; a = 12; b = 36;
#1; a = 12; b = 37;
#1; a = 12; b = 38;
#1; a = 12; b = 39;
#1; a = 13; b = 0;
#1; a = 13; b = 1;
#1; a = 13; b = 2;
#1; a = 13; b = 3;
#1; a = 13; b = 4;
#1; a = 13; b = 5;
#1; a = 13; b = 6;
#1; a = 13; b = 7;
#1; a = 13; b = 8;
#1; a = 13; b = 9;
#1; a = 13; b = 10;
#1; a = 13; b = 11;
#1; a = 13; b = 12;
#1; a = 13; b = 13;
#1; a = 13; b = 14;
#1; a = 13; b = 15;
#1; a = 13; b = 16;
#1; a = 13; b = 17;
#1; a = 13; b = 18;
#1; a = 13; b = 19;
#1; a = 13; b = 20;
#1; a = 13; b = 21;
#1; a = 13; b = 22;
#1; a = 13; b = 23;
#1; a = 13; b = 24;
#1; a = 13; b = 25;
#1; a = 13; b = 26;
#1; a = 13; b = 27;
#1; a = 13; b = 28;
#1; a = 13; b = 29;
#1; a = 13; b = 30;
#1; a = 13; b = 31;
#1; a = 13; b = 32;
#1; a = 13; b = 33;
#1; a = 13; b = 34;
#1; a = 13; b = 35;
#1; a = 13; b = 36;
#1; a = 13; b = 37;
#1; a = 13; b = 38;
#1; a = 13; b = 39;
#1; a = 14; b = 0;
#1; a = 14; b = 1;
#1; a = 14; b = 2;
#1; a = 14; b = 3;
#1; a = 14; b = 4;
#1; a = 14; b = 5;
#1; a = 14; b = 6;
#1; a = 14; b = 7;
#1; a = 14; b = 8;
#1; a = 14; b = 9;
#1; a = 14; b = 10;
#1; a = 14; b = 11;
#1; a = 14; b = 12;
#1; a = 14; b = 13;
#1; a = 14; b = 14;
#1; a = 14; b = 15;
#1; a = 14; b = 16;
#1; a = 14; b = 17;
#1; a = 14; b = 18;
#1; a = 14; b = 19;
#1; a = 14; b = 20;
#1; a = 14; b = 21;
#1; a = 14; b = 22;
#1; a = 14; b = 23;
#1; a = 14; b = 24;
#1; a = 14; b = 25;
#1; a = 14; b = 26;
#1; a = 14; b = 27;
#1; a = 14; b = 28;
#1; a = 14; b = 29;
#1; a = 14; b = 30;
#1; a = 14; b = 31;
#1; a = 14; b = 32;
#1; a = 14; b = 33;
#1; a = 14; b = 34;
#1; a = 14; b = 35;
#1; a = 14; b = 36;
#1; a = 14; b = 37;
#1; a = 14; b = 38;
#1; a = 14; b = 39;
#1; a = 15; b = 0;
#1; a = 15; b = 1;
#1; a = 15; b = 2;
#1; a = 15; b = 3;
#1; a = 15; b = 4;
#1; a = 15; b = 5;
#1; a = 15; b = 6;
#1; a = 15; b = 7;
#1; a = 15; b = 8;
#1; a = 15; b = 9;
#1; a = 15; b = 10;
#1; a = 15; b = 11;
#1; a = 15; b = 12;
#1; a = 15; b = 13;
#1; a = 15; b = 14;
#1; a = 15; b = 15;
#1; a = 15; b = 16;
#1; a = 15; b = 17;
#1; a = 15; b = 18;
#1; a = 15; b = 19;
#1; a = 15; b = 20;
#1; a = 15; b = 21;
#1; a = 15; b = 22;
#1; a = 15; b = 23;
#1; a = 15; b = 24;
#1; a = 15; b = 25;
#1; a = 15; b = 26;
#1; a = 15; b = 27;
#1; a = 15; b = 28;
#1; a = 15; b = 29;
#1; a = 15; b = 30;
#1; a = 15; b = 31;
#1; a = 15; b = 32;
#1; a = 15; b = 33;
#1; a = 15; b = 34;
#1; a = 15; b = 35;
#1; a = 15; b = 36;
#1; a = 15; b = 37;
#1; a = 15; b = 38;
#1; a = 15; b = 39;

        #10; $finish;
    end
endmodule
