`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05.12.2024 13:19:09
// Design Name: 
// Module Name: CharacterIdEncoderTest
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module CharacterIdEncoderTest(

    );
    
    wire [7:0] character_id;
    reg [7:0] input_id;
    reg clock;
    
    CharacterIdEncoder characterIdEncoder(character_id,input_id,1,clock);
    
    initial begin
        input_id = 0;
        clock = 0;
        #1; input_id = 0;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 1;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 2;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 3;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 4;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 5;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 6;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 7;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 8;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 9;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 10;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 11;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 12;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 13;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 14;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 15;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 16;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 17;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 18;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 19;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 20;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 21;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 22;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 23;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 24;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 25;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 26;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 27;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 28;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 29;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 30;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 31;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 32;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 33;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 34;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 35;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 36;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 37;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 38;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 39;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 40;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 41;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 42;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 43;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 44;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 45;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 46;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 47;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 48;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 49;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 50;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 51;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 52;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 53;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 54;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 55;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 56;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 57;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 58;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 59;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 60;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 61;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 62;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 63;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 64;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 65;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 66;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 67;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 68;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 69;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 70;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 71;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 72;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 73;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 74;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 75;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 76;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 77;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 78;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 79;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 80;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 81;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 82;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 83;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 84;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 85;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 86;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 87;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 88;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 89;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 90;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 91;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 92;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 93;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 94;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 95;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 96;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 97;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 98;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 99;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 100;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 101;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 102;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 103;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 104;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 105;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 106;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 107;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 108;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 109;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 110;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 111;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 112;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 113;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 114;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 115;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 116;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 117;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 118;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 119;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 120;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 121;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 122;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 123;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 124;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 125;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 126;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 127;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 128;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 129;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 130;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 131;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 132;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 133;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 134;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 135;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 136;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 137;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 138;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 139;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 140;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 141;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 142;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 143;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 144;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 145;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 146;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 147;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 148;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 149;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 150;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 151;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 152;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 153;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 154;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 155;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 156;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 157;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 158;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 159;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 160;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 161;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 162;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 163;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 164;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 165;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 166;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 167;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 168;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 169;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 170;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 171;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 172;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 173;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 174;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 175;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 176;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 177;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 178;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 179;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 180;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 181;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 182;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 183;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 184;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 185;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 186;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 187;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 188;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 189;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 190;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 191;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 192;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 193;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 194;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 195;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 196;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 197;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 198;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 199;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 200;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 201;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 202;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 203;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 204;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 205;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 206;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 207;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 208;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 209;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 210;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 211;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 212;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 213;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 214;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 215;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 216;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 217;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 218;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 219;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 220;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 221;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 222;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 223;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 224;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 225;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 226;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 227;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 228;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 229;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 230;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 231;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 232;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 233;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 234;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 235;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 236;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 237;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 238;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 239;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 240;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 241;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 242;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 243;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 244;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 245;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 246;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 247;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 248;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 249;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 250;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 251;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 252;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 253;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 254;
        #1; clock = 1;
        #1; clock = 0;
        #1; input_id = 255;
        #1; clock = 1;
        #1; clock = 0;

    end
    
endmodule
